module vlang_page_parser

pub fn parse_html(html_string string) string {
	return html_string
}
